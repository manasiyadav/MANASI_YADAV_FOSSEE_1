* C:\Users\admin\eSim-Workspace\priencoder\priencoder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/15/21 19:51:08

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ priencoder		
U2  Net-_R1-Pad2_ Net-_R2-Pad2_ Net-_R3-Pad2_ Net-_R4-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ adc_bridge_4		
U3  Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_R7-Pad2_ Net-_R6-Pad2_ Net-_R5-Pad2_ dac_bridge_3		
R7  Net-_R1-Pad1_ Net-_R7-Pad2_ 100k		
R4  Net-_R1-Pad1_ Net-_R4-Pad2_ 100k		
v4  Net-_R4-Pad2_ Net-_R1-Pad1_ pulse		
R3  Net-_R1-Pad1_ Net-_R3-Pad2_ 100k		
v3  Net-_R3-Pad2_ Net-_R1-Pad1_ pulse		
R2  Net-_R1-Pad1_ Net-_R2-Pad2_ 100k		
v2  Net-_R2-Pad2_ Net-_R1-Pad1_ pulse		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 100k		
v1  Net-_R1-Pad2_ Net-_R1-Pad1_ pulse		
R5  Net-_R1-Pad1_ Net-_R5-Pad2_ 100k		
R6  Net-_R1-Pad1_ Net-_R6-Pad2_ 100k		

.end
